package ula_package is

	type ULA_OPERATION is (ADD);

end package;